class Integer {
    int value;
    long hash() {
        return self.value;
    }
}

class Long {
    long value;
    long hash() {
        return self.value;
    }
}

class Short {
    short value;
    long hash() {
        return self.value;
    }
}

class Char {
    char value;
    long hash() {
        return self.value;
    }
}

class Float {
    float value;
    long hash() {
        return self.value;
    }
}

class Double {
    double value;
    long hash() {
        return self.value;
    }
}
