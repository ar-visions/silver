include stdlib;

class Super {
    void super_only(int test) {
        printf("super only");
    }
    void method(int arg, int arg2) {
        printf("original function");
    }
}